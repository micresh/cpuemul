module ALU_tb;
	
	reg [7:0] A = 8'b00000000;
	reg [7:0]

endmodule;
